magic
tech sky130A
timestamp 1616446594
<< nwell >>
rect 472 77 600 413
<< nmos >>
rect 530 -95 545 5
<< pmos >>
rect 530 95 545 395
<< ndiff >>
rect 490 -10 530 5
rect 490 -27 495 -10
rect 512 -27 530 -10
rect 490 -63 530 -27
rect 490 -80 495 -63
rect 512 -80 530 -63
rect 490 -95 530 -80
rect 545 -10 582 5
rect 545 -27 558 -10
rect 575 -27 582 -10
rect 545 -63 582 -27
rect 545 -80 558 -63
rect 575 -80 582 -63
rect 545 -95 582 -80
<< pdiff >>
rect 490 380 530 395
rect 490 363 495 380
rect 512 363 530 380
rect 490 257 530 363
rect 490 240 495 257
rect 512 240 530 257
rect 490 127 530 240
rect 490 110 495 127
rect 512 110 530 127
rect 490 95 530 110
rect 545 380 582 395
rect 545 363 558 380
rect 575 363 582 380
rect 545 257 582 363
rect 545 240 558 257
rect 575 240 582 257
rect 545 127 582 240
rect 545 110 558 127
rect 575 110 582 127
rect 545 95 582 110
<< ndiffc >>
rect 495 -27 512 -10
rect 495 -80 512 -63
rect 558 -27 575 -10
rect 558 -80 575 -63
<< pdiffc >>
rect 495 363 512 380
rect 495 240 512 257
rect 495 110 512 127
rect 558 363 575 380
rect 558 240 575 257
rect 558 110 575 127
<< poly >>
rect 530 395 545 417
rect 416 56 453 67
rect 416 39 426 56
rect 443 55 453 56
rect 530 55 545 95
rect 443 39 545 55
rect 416 38 545 39
rect 416 30 453 38
rect 530 5 545 38
rect 530 -125 545 -95
<< polycont >>
rect 426 39 443 56
<< locali >>
rect 508 460 530 477
rect 547 460 566 477
rect 495 380 512 460
rect 495 257 512 363
rect 495 127 512 240
rect 495 100 512 110
rect 558 380 575 390
rect 558 257 575 363
rect 558 127 575 240
rect 416 56 453 67
rect 416 39 426 56
rect 443 39 453 56
rect 416 30 453 39
rect 558 55 575 110
rect 649 55 686 65
rect 558 38 686 55
rect 495 -10 512 0
rect 495 -63 512 -27
rect 495 -180 512 -80
rect 558 -10 575 38
rect 649 28 686 38
rect 558 -63 575 -27
rect 558 -90 575 -80
rect 507 -197 529 -180
rect 546 -197 567 -180
<< viali >>
rect 491 460 508 477
rect 530 460 547 477
rect 566 460 583 477
rect 490 -197 507 -180
rect 529 -197 546 -180
rect 567 -197 584 -180
<< metal1 >>
rect 480 477 590 485
rect 480 460 491 477
rect 508 460 530 477
rect 547 460 566 477
rect 583 460 590 477
rect 480 450 590 460
rect 480 -180 590 -170
rect 480 -197 490 -180
rect 507 -197 529 -180
rect 546 -197 567 -180
rect 584 -197 590 -180
rect 480 -205 590 -197
<< labels >>
flabel polycont 426 39 443 56 0 FreeSans 80 0 0 0 in
flabel viali 529 -197 546 -180 0 FreeSans 80 0 0 0 vgnd
flabel locali 660 38 677 55 0 FreeSans 80 0 0 0 out
flabel viali 530 460 547 477 0 FreeSans 80 0 0 0 vdd
flabel space 558 -162 575 -145 0 FreeSans 80 0 0 0 pbulk
flabel space 583 397 600 414 0 FreeSans 80 0 0 0 nbulk
<< end >>
